module not_gate (a,b);
integer a;

input a
input b

assign b = ~a

endmodule



